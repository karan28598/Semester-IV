*Clipper Circuit without bias
Vin 1 0 sin(5V 0V 1khz)
R1 2 1 1.1k
Diode 0 2 D2
.model D2 D
.tran 0 5ms
.probe
.end