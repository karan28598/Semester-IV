*Full Wave Rectifier LC Filter
Vin 5 0 sin(0 230V 50Hz)
r1 1 5 1k
l1 1 0 0.5h
l2 2 0 0.5h
l3 3 0 0.5h
k1 l1 l2 0.999
k2 l1 l3 0.999
k3 l2 l3 0.999
d1 2 4 diode
d2 3 4 diode
l4 4 6 1
c 4 0 10uf
r2 6 0 470
.model diode d
.tran 0 50ms
.probe
.end