*Full Wave Rectifier PI Filter
Vin 6 0 sin(0 230V 50Hz)
r1 6 1 0.3
l1 1 0 0.5h
l2 2 0 0.5h
l3 0 3 0.5h
k12 l1 l2 0.999
k23 l2 l3 0.999
k31 l3 l1 0.999
d1 2 4 diode
d2 3 4 diode
R 5 0 0.5k
l 4 5 1000mh
c1 4 0 10u
c2 5 0 10u
.model diode d
.tran 0ms 80ms
.probe
.end