*Zener Diode Forward Bias
Vin 1 0 10Vdc
r 1 2 1k
d 0 2 zener
.model zenerd(bv=2v)
.dc Vin -10 10 0.5v
.probe
.end