*BJT Characteristics Voltage Divider
vbb 1 0 0v
vcc 3 0 0v
r1 1 2 12k
r2 1 0 4.5k
rc 5 2 470
re 6 0 70
q 5 1 6 BJT
.model BJT npm(ls=10E-16,Bf=220,Va=100V,CJe=5pf)
.Dc vbb 0 10v .1v vcc 0 3v 1v
.probe
.end